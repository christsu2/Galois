/* Bleen Systems, Inc. Confidential Information */
/* Copyright (C) 2003 Baleen Systems, Inc. */

/* $Header: L:\\src/lightning2/rtl/ECC/rsROM.v,v 1.1 2003/05/27 17:34:54 JEROME Exp $ */
/*---------------------------------------------------------------------------*
 * Author            : Hon-Ming Li
 * Created on        : Wed March 19 10:34:28 PST 2003
 * Last checked in by: $Author: JEROME $
 * Last checked in on: $Date: 2003/05/27 17:34:54 $
 *
 *---------------------------------------------------------------------------*/
/*
 * $Log: rsROM.v,v $
 * Revision 1.1  2003/05/27 17:34:54  JEROME
 * *** empty log message ***
 *
 * Revision 1.3  2003/04/29 00:50:05  mingl
 * new code with results in "absolute byte location"
 *
 * Revision 1.2  2003/03/19 18:41:03  mingl
 * add CVS header, change initial value of state machine (from 8'hxx to 8'h00)
 *
 *
 */

module rsROM(i, q);
input [8:0] i;
output[7:0] q;

reg[7:0] q;

always @(i)


case(i)
//invert table

   0: q =   1;
   1: q =   1;
   2: q = 142;
   3: q = 244;
   4: q =  71;
   5: q = 167;
   6: q = 122;
   7: q = 186;
   8: q = 173;
   9: q = 157;
  10: q = 221;
  11: q = 152;
  12: q =  61;
  13: q = 170;
  14: q =  93;
  15: q = 150;
  16: q = 216;
  17: q = 114;
  18: q = 192;
  19: q =  88;
  20: q = 224;
  21: q =  62;
  22: q =  76;
  23: q = 102;
  24: q = 144;
  25: q = 222;
  26: q =  85;
  27: q = 128;
  28: q = 160;
  29: q = 131;
  30: q =  75;
  31: q =  42;
  32: q = 108;
  33: q = 237;
  34: q =  57;
  35: q =  81;
  36: q =  96;
  37: q =  86;
  38: q =  44;
  39: q = 138;
  40: q = 112;
  41: q = 208;
  42: q =  31;
  43: q =  74;
  44: q =  38;
  45: q = 139;
  46: q =  51;
  47: q = 110;
  48: q =  72;
  49: q = 137;
  50: q = 111;
  51: q =  46;
  52: q = 164;
  53: q = 195;
  54: q =  64;
  55: q =  94;
  56: q =  80;
  57: q =  34;
  58: q = 207;
  59: q = 169;
  60: q = 171;
  61: q =  12;
  62: q =  21;
  63: q = 225;
  64: q =  54;
  65: q =  95;
  66: q = 248;
  67: q = 213;
  68: q = 146;
  69: q =  78;
  70: q = 166;
  71: q =   4;
  72: q =  48;
  73: q = 136;
  74: q =  43;
  75: q =  30;
  76: q =  22;
  77: q = 103;
  78: q =  69;
  79: q = 147;
  80: q =  56;
  81: q =  35;
  82: q = 104;
  83: q = 140;
  84: q = 129;
  85: q =  26;
  86: q =  37;
  87: q =  97;
  88: q =  19;
  89: q = 193;
  90: q = 203;
  91: q =  99;
  92: q = 151;
  93: q =  14;
  94: q =  55;
  95: q =  65;
  96: q =  36;
  97: q =  87;
  98: q = 202;
  99: q =  91;
 100: q = 185;
 101: q = 196;
 102: q =  23;
 103: q =  77;
 104: q =  82;
 105: q = 141;
 106: q = 239;
 107: q = 179;
 108: q =  32;
 109: q = 236;
 110: q =  47;
 111: q =  50;
 112: q =  40;
 113: q = 209;
 114: q =  17;
 115: q = 217;
 116: q = 233;
 117: q = 251;
 118: q = 218;
 119: q = 121;
 120: q = 219;
 121: q = 119;
 122: q =   6;
 123: q = 187;
 124: q = 132;
 125: q = 205;
 126: q = 254;
 127: q = 252;
 128: q =  27;
 129: q =  84;
 130: q = 161;
 131: q =  29;
 132: q = 124;
 133: q = 204;
 134: q = 228;
 135: q = 176;
 136: q =  73;
 137: q =  49;
 138: q =  39;
 139: q =  45;
 140: q =  83;
 141: q = 105;
 142: q =   2;
 143: q = 245;
 144: q =  24;
 145: q = 223;
 146: q =  68;
 147: q =  79;
 148: q = 155;
 149: q = 188;
 150: q =  15;
 151: q =  92;
 152: q =  11;
 153: q = 220;
 154: q = 189;
 155: q = 148;
 156: q = 172;
 157: q =   9;
 158: q = 199;
 159: q = 162;
 160: q =  28;
 161: q = 130;
 162: q = 159;
 163: q = 198;
 164: q =  52;
 165: q = 194;
 166: q =  70;
 167: q =   5;
 168: q = 206;
 169: q =  59;
 170: q =  13;
 171: q =  60;
 172: q = 156;
 173: q =   8;
 174: q = 190;
 175: q = 183;
 176: q = 135;
 177: q = 229;
 178: q = 238;
 179: q = 107;
 180: q = 235;
 181: q = 242;
 182: q = 191;
 183: q = 175;
 184: q = 197;
 185: q = 100;
 186: q =   7;
 187: q = 123;
 188: q = 149;
 189: q = 154;
 190: q = 174;
 191: q = 182;
 192: q =  18;
 193: q =  89;
 194: q = 165;
 195: q =  53;
 196: q = 101;
 197: q = 184;
 198: q = 163;
 199: q = 158;
 200: q = 210;
 201: q = 247;
 202: q =  98;
 203: q =  90;
 204: q = 133;
 205: q = 125;
 206: q = 168;
 207: q =  58;
 208: q =  41;
 209: q = 113;
 210: q = 200;
 211: q = 246;
 212: q = 249;
 213: q =  67;
 214: q = 215;
 215: q = 214;
 216: q =  16;
 217: q = 115;
 218: q = 118;
 219: q = 120;
 220: q = 153;
 221: q =  10;
 222: q =  25;
 223: q = 145;
 224: q =  20;
 225: q =  63;
 226: q = 230;
 227: q = 240;
 228: q = 134;
 229: q = 177;
 230: q = 226;
 231: q = 241;
 232: q = 250;
 233: q = 116;
 234: q = 243;
 235: q = 180;
 236: q = 109;
 237: q =  33;
 238: q = 178;
 239: q = 106;
 240: q = 227;
 241: q = 231;
 242: q = 181;
 243: q = 234;
 244: q =   3;
 245: q = 143;
 246: q = 211;
 247: q = 201;
 248: q =  66;
 249: q = 212;
 250: q = 232;
 251: q = 117;
 252: q = 127;
 253: q = 255;
 254: q = 126;
 255: q = 253;

//Antilog Table

 256: q = 255;
 257: q =   0;
 258: q =   1;
 259: q =  25;
 260: q =   2;
 261: q =  50;
 262: q =  26;
 263: q = 198;
 264: q =   3;
 265: q = 223;
 266: q =  51;
 267: q = 238;
 268: q =  27;
 269: q = 104;
 270: q = 199;
 271: q =  75;
 272: q =   4;
 273: q = 100;
 274: q = 224;
 275: q =  14;
 276: q =  52;
 277: q = 141;
 278: q = 239;
 279: q = 129;
 280: q =  28;
 281: q = 193;
 282: q = 105;
 283: q = 248;
 284: q = 200;
 285: q =   8;
 286: q =  76;
 287: q = 113;
 288: q =   5;
 289: q = 138;
 290: q = 101;
 291: q =  47;
 292: q = 225;
 293: q =  36;
 294: q =  15;
 295: q =  33;
 296: q =  53;
 297: q = 147;
 298: q = 142;
 299: q = 218;
 300: q = 240;
 301: q =  18;
 302: q = 130;
 303: q =  69;
 304: q =  29;
 305: q = 181;
 306: q = 194;
 307: q = 125;
 308: q = 106;
 309: q =  39;
 310: q = 249;
 311: q = 185;
 312: q = 201;
 313: q = 154;
 314: q =   9;
 315: q = 120;
 316: q =  77;
 317: q = 228;
 318: q = 114;
 319: q = 166;
 320: q =   6;
 321: q = 191;
 322: q = 139;
 323: q =  98;
 324: q = 102;
 325: q = 221;
 326: q =  48;
 327: q = 253;
 328: q = 226;
 329: q = 152;
 330: q =  37;
 331: q = 179;
 332: q =  16;
 333: q = 145;
 334: q =  34;
 335: q = 136;
 336: q =  54;
 337: q = 208;
 338: q = 148;
 339: q = 206;
 340: q = 143;
 341: q = 150;
 342: q = 219;
 343: q = 189;
 344: q = 241;
 345: q = 210;
 346: q =  19;
 347: q =  92;
 348: q = 131;
 349: q =  56;
 350: q =  70;
 351: q =  64;
 352: q =  30;
 353: q =  66;
 354: q = 182;
 355: q = 163;
 356: q = 195;
 357: q =  72;
 358: q = 126;
 359: q = 110;
 360: q = 107;
 361: q =  58;
 362: q =  40;
 363: q =  84;
 364: q = 250;
 365: q = 133;
 366: q = 186;
 367: q =  61;
 368: q = 202;
 369: q =  94;
 370: q = 155;
 371: q = 159;
 372: q =  10;
 373: q =  21;
 374: q = 121;
 375: q =  43;
 376: q =  78;
 377: q = 212;
 378: q = 229;
 379: q = 172;
 380: q = 115;
 381: q = 243;
 382: q = 167;
 383: q =  87;
 384: q =   7;
 385: q = 112;
 386: q = 192;
 387: q = 247;
 388: q = 140;
 389: q = 128;
 390: q =  99;
 391: q =  13;
 392: q = 103;
 393: q =  74;
 394: q = 222;
 395: q = 237;
 396: q =  49;
 397: q = 197;
 398: q = 254;
 399: q =  24;
 400: q = 227;
 401: q = 165;
 402: q = 153;
 403: q = 119;
 404: q =  38;
 405: q = 184;
 406: q = 180;
 407: q = 124;
 408: q =  17;
 409: q =  68;
 410: q = 146;
 411: q = 217;
 412: q =  35;
 413: q =  32;
 414: q = 137;
 415: q =  46;
 416: q =  55;
 417: q =  63;
 418: q = 209;
 419: q =  91;
 420: q = 149;
 421: q = 188;
 422: q = 207;
 423: q = 205;
 424: q = 144;
 425: q = 135;
 426: q = 151;
 427: q = 178;
 428: q = 220;
 429: q = 252;
 430: q = 190;
 431: q =  97;
 432: q = 242;
 433: q =  86;
 434: q = 211;
 435: q = 171;
 436: q =  20;
 437: q =  42;
 438: q =  93;
 439: q = 158;
 440: q = 132;
 441: q =  60;
 442: q =  57;
 443: q =  83;
 444: q =  71;
 445: q = 109;
 446: q =  65;
 447: q = 162;
 448: q =  31;
 449: q =  45;
 450: q =  67;
 451: q = 216;
 452: q = 183;
 453: q = 123;
 454: q = 164;
 455: q = 118;
 456: q = 196;
 457: q =  23;
 458: q =  73;
 459: q = 236;
 460: q = 127;
 461: q =  12;
 462: q = 111;
 463: q = 246;
 464: q = 108;
 465: q = 161;
 466: q =  59;
 467: q =  82;
 468: q =  41;
 469: q = 157;
 470: q =  85;
 471: q = 170;
 472: q = 251;
 473: q =  96;
 474: q = 134;
 475: q = 177;
 476: q = 187;
 477: q = 204;
 478: q =  62;
 479: q =  90;
 480: q = 203;
 481: q =  89;
 482: q =  95;
 483: q = 176;
 484: q = 156;
 485: q = 169;
 486: q = 160;
 487: q =  81;
 488: q =  11;
 489: q = 245;
 490: q =  22;
 491: q = 235;
 492: q = 122;
 493: q = 117;
 494: q =  44;
 495: q = 215;
 496: q =  79;
 497: q = 174;
 498: q = 213;
 499: q = 233;
 500: q = 230;
 501: q = 231;
 502: q = 173;
 503: q = 232;
 504: q = 116;
 505: q = 214;
 506: q = 244;
 507: q = 234;
 508: q = 168;
 509: q =  80;
 510: q =  88;
 511: q = 175;

endcase
endmodule
