module rsROM(i, q, clk);
input [8:0] i;
input       clk;
output[7:0] q;

reg[7:0] x, q;

always @(posedge clk)
     q <= #1 x;         
	
always @(i)
case(i)
//invert table

   0: x =   1;
   1: x =   1;
   2: x = 142;
   3: x = 244;
   4: x =  71;
   5: x = 167;
   6: x = 122;
   7: x = 186;
   8: x = 173;
   9: x = 157;
  10: x = 221;
  11: x = 152;
  12: x =  61;
  13: x = 170;
  14: x =  93;
  15: x = 150;
  16: x = 216;
  17: x = 114;
  18: x = 192;
  19: x =  88;
  20: x = 224;
  21: x =  62;
  22: x =  76;
  23: x = 102;
  24: x = 144;
  25: x = 222;
  26: x =  85;
  27: x = 128;
  28: x = 160;
  29: x = 131;
  30: x =  75;
  31: x =  42;
  32: x = 108;
  33: x = 237;
  34: x =  57;
  35: x =  81;
  36: x =  96;
  37: x =  86;
  38: x =  44;
  39: x = 138;
  40: x = 112;
  41: x = 208;
  42: x =  31;
  43: x =  74;
  44: x =  38;
  45: x = 139;
  46: x =  51;
  47: x = 110;
  48: x =  72;
  49: x = 137;
  50: x = 111;
  51: x =  46;
  52: x = 164;
  53: x = 195;
  54: x =  64;
  55: x =  94;
  56: x =  80;
  57: x =  34;
  58: x = 207;
  59: x = 169;
  60: x = 171;
  61: x =  12;
  62: x =  21;
  63: x = 225;
  64: x =  54;
  65: x =  95;
  66: x = 248;
  67: x = 213;
  68: x = 146;
  69: x =  78;
  70: x = 166;
  71: x =   4;
  72: x =  48;
  73: x = 136;
  74: x =  43;
  75: x =  30;
  76: x =  22;
  77: x = 103;
  78: x =  69;
  79: x = 147;
  80: x =  56;
  81: x =  35;
  82: x = 104;
  83: x = 140;
  84: x = 129;
  85: x =  26;
  86: x =  37;
  87: x =  97;
  88: x =  19;
  89: x = 193;
  90: x = 203;
  91: x =  99;
  92: x = 151;
  93: x =  14;
  94: x =  55;
  95: x =  65;
  96: x =  36;
  97: x =  87;
  98: x = 202;
  99: x =  91;
 100: x = 185;
 101: x = 196;
 102: x =  23;
 103: x =  77;
 104: x =  82;
 105: x = 141;
 106: x = 239;
 107: x = 179;
 108: x =  32;
 109: x = 236;
 110: x =  47;
 111: x =  50;
 112: x =  40;
 113: x = 209;
 114: x =  17;
 115: x = 217;
 116: x = 233;
 117: x = 251;
 118: x = 218;
 119: x = 121;
 120: x = 219;
 121: x = 119;
 122: x =   6;
 123: x = 187;
 124: x = 132;
 125: x = 205;
 126: x = 254;
 127: x = 252;
 128: x =  27;
 129: x =  84;
 130: x = 161;
 131: x =  29;
 132: x = 124;
 133: x = 204;
 134: x = 228;
 135: x = 176;
 136: x =  73;
 137: x =  49;
 138: x =  39;
 139: x =  45;
 140: x =  83;
 141: x = 105;
 142: x =   2;
 143: x = 245;
 144: x =  24;
 145: x = 223;
 146: x =  68;
 147: x =  79;
 148: x = 155;
 149: x = 188;
 150: x =  15;
 151: x =  92;
 152: x =  11;
 153: x = 220;
 154: x = 189;
 155: x = 148;
 156: x = 172;
 157: x =   9;
 158: x = 199;
 159: x = 162;
 160: x =  28;
 161: x = 130;
 162: x = 159;
 163: x = 198;
 164: x =  52;
 165: x = 194;
 166: x =  70;
 167: x =   5;
 168: x = 206;
 169: x =  59;
 170: x =  13;
 171: x =  60;
 172: x = 156;
 173: x =   8;
 174: x = 190;
 175: x = 183;
 176: x = 135;
 177: x = 229;
 178: x = 238;
 179: x = 107;
 180: x = 235;
 181: x = 242;
 182: x = 191;
 183: x = 175;
 184: x = 197;
 185: x = 100;
 186: x =   7;
 187: x = 123;
 188: x = 149;
 189: x = 154;
 190: x = 174;
 191: x = 182;
 192: x =  18;
 193: x =  89;
 194: x = 165;
 195: x =  53;
 196: x = 101;
 197: x = 184;
 198: x = 163;
 199: x = 158;
 200: x = 210;
 201: x = 247;
 202: x =  98;
 203: x =  90;
 204: x = 133;
 205: x = 125;
 206: x = 168;
 207: x =  58;
 208: x =  41;
 209: x = 113;
 210: x = 200;
 211: x = 246;
 212: x = 249;
 213: x =  67;
 214: x = 215;
 215: x = 214;
 216: x =  16;
 217: x = 115;
 218: x = 118;
 219: x = 120;
 220: x = 153;
 221: x =  10;
 222: x =  25;
 223: x = 145;
 224: x =  20;
 225: x =  63;
 226: x = 230;
 227: x = 240;
 228: x = 134;
 229: x = 177;
 230: x = 226;
 231: x = 241;
 232: x = 250;
 233: x = 116;
 234: x = 243;
 235: x = 180;
 236: x = 109;
 237: x =  33;
 238: x = 178;
 239: x = 106;
 240: x = 227;
 241: x = 231;
 242: x = 181;
 243: x = 234;
 244: x =   3;
 245: x = 143;
 246: x = 211;
 247: x = 201;
 248: x =  66;
 249: x = 212;
 250: x = 232;
 251: x = 117;
 252: x = 127;
 253: x = 255;
 254: x = 126;
 255: x = 253;

//Antilog Table

 256: x = 255;
 257: x =   0;
 258: x =   1;
 259: x =  25;
 260: x =   2;
 261: x =  50;
 262: x =  26;
 263: x = 198;
 264: x =   3;
 265: x = 223;
 266: x =  51;
 267: x = 238;
 268: x =  27;
 269: x = 104;
 270: x = 199;
 271: x =  75;
 272: x =   4;
 273: x = 100;
 274: x = 224;
 275: x =  14;
 276: x =  52;
 277: x = 141;
 278: x = 239;
 279: x = 129;
 280: x =  28;
 281: x = 193;
 282: x = 105;
 283: x = 248;
 284: x = 200;
 285: x =   8;
 286: x =  76;
 287: x = 113;
 288: x =   5;
 289: x = 138;
 290: x = 101;
 291: x =  47;
 292: x = 225;
 293: x =  36;
 294: x =  15;
 295: x =  33;
 296: x =  53;
 297: x = 147;
 298: x = 142;
 299: x = 218;
 300: x = 240;
 301: x =  18;
 302: x = 130;
 303: x =  69;
 304: x =  29;
 305: x = 181;
 306: x = 194;
 307: x = 125;
 308: x = 106;
 309: x =  39;
 310: x = 249;
 311: x = 185;
 312: x = 201;
 313: x = 154;
 314: x =   9;
 315: x = 120;
 316: x =  77;
 317: x = 228;
 318: x = 114;
 319: x = 166;
 320: x =   6;
 321: x = 191;
 322: x = 139;
 323: x =  98;
 324: x = 102;
 325: x = 221;
 326: x =  48;
 327: x = 253;
 328: x = 226;
 329: x = 152;
 330: x =  37;
 331: x = 179;
 332: x =  16;
 333: x = 145;
 334: x =  34;
 335: x = 136;
 336: x =  54;
 337: x = 208;
 338: x = 148;
 339: x = 206;
 340: x = 143;
 341: x = 150;
 342: x = 219;
 343: x = 189;
 344: x = 241;
 345: x = 210;
 346: x =  19;
 347: x =  92;
 348: x = 131;
 349: x =  56;
 350: x =  70;
 351: x =  64;
 352: x =  30;
 353: x =  66;
 354: x = 182;
 355: x = 163;
 356: x = 195;
 357: x =  72;
 358: x = 126;
 359: x = 110;
 360: x = 107;
 361: x =  58;
 362: x =  40;
 363: x =  84;
 364: x = 250;
 365: x = 133;
 366: x = 186;
 367: x =  61;
 368: x = 202;
 369: x =  94;
 370: x = 155;
 371: x = 159;
 372: x =  10;
 373: x =  21;
 374: x = 121;
 375: x =  43;
 376: x =  78;
 377: x = 212;
 378: x = 229;
 379: x = 172;
 380: x = 115;
 381: x = 243;
 382: x = 167;
 383: x =  87;
 384: x =   7;
 385: x = 112;
 386: x = 192;
 387: x = 247;
 388: x = 140;
 389: x = 128;
 390: x =  99;
 391: x =  13;
 392: x = 103;
 393: x =  74;
 394: x = 222;
 395: x = 237;
 396: x =  49;
 397: x = 197;
 398: x = 254;
 399: x =  24;
 400: x = 227;
 401: x = 165;
 402: x = 153;
 403: x = 119;
 404: x =  38;
 405: x = 184;
 406: x = 180;
 407: x = 124;
 408: x =  17;
 409: x =  68;
 410: x = 146;
 411: x = 217;
 412: x =  35;
 413: x =  32;
 414: x = 137;
 415: x =  46;
 416: x =  55;
 417: x =  63;
 418: x = 209;
 419: x =  91;
 420: x = 149;
 421: x = 188;
 422: x = 207;
 423: x = 205;
 424: x = 144;
 425: x = 135;
 426: x = 151;
 427: x = 178;
 428: x = 220;
 429: x = 252;
 430: x = 190;
 431: x =  97;
 432: x = 242;
 433: x =  86;
 434: x = 211;
 435: x = 171;
 436: x =  20;
 437: x =  42;
 438: x =  93;
 439: x = 158;
 440: x = 132;
 441: x =  60;
 442: x =  57;
 443: x =  83;
 444: x =  71;
 445: x = 109;
 446: x =  65;
 447: x = 162;
 448: x =  31;
 449: x =  45;
 450: x =  67;
 451: x = 216;
 452: x = 183;
 453: x = 123;
 454: x = 164;
 455: x = 118;
 456: x = 196;
 457: x =  23;
 458: x =  73;
 459: x = 236;
 460: x = 127;
 461: x =  12;
 462: x = 111;
 463: x = 246;
 464: x = 108;
 465: x = 161;
 466: x =  59;
 467: x =  82;
 468: x =  41;
 469: x = 157;
 470: x =  85;
 471: x = 170;
 472: x = 251;
 473: x =  96;
 474: x = 134;
 475: x = 177;
 476: x = 187;
 477: x = 204;
 478: x =  62;
 479: x =  90;
 480: x = 203;
 481: x =  89;
 482: x =  95;
 483: x = 176;
 484: x = 156;
 485: x = 169;
 486: x = 160;
 487: x =  81;
 488: x =  11;
 489: x = 245;
 490: x =  22;
 491: x = 235;
 492: x = 122;
 493: x = 117;
 494: x =  44;
 495: x = 215;
 496: x =  79;
 497: x = 174;
 498: x = 213;
 499: x = 233;
 500: x = 230;
 501: x = 231;
 502: x = 173;
 503: x = 232;
 504: x = 116;
 505: x = 214;
 506: x = 244;
 507: x = 234;
 508: x = 168;
 509: x =  80;
 510: x =  88;
 511: x = 175;

endcase
endmodule
